module tfgrid

//logic needs to be here to fetch basic info from TFGrid DB

struct Explorer{

	ipaddr: []string

}


fn explorer_new ()? Explorer{

	mut explorer := Explorer{}

	//now add the ipaddresses in code which explorers can be reached


}