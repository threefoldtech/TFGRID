module tfgrid

pub struct PublicIP {
pub mut:
	ip string
}

pub struct PublicIPResult {
pub mut:
	ip string
}
