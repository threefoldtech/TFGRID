
module tfgrid

//as registered on the TFGrid DB
struct TFGridEntity{

}

struct TFGridTwin{

}

struct TFGridNode{

}

struct TFGridFarmer{

}