
module tfgrid

//as registered on the TFGrid DB
//need the data models here
struct TFGridEntity{

}

struct TFGridTwin{

}

struct TFGridNode{

}

struct TFGridFarmer{

}