module tfgrid

struct MyTwin {}

fn (mut grid MyTwin) init() ? {
}
